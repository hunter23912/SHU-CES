`default_nettype none

/* verilator lint_off BLKSEQ */

`include "Lock.v"

module tb_Lock ();
  reg clk_tb;//ʱ���ź�
  reg rst_n_tb;//��λ�ź�
  reg modeSettingWire_tb;//��������ģʽ
  reg inputNextSignal_tb;//������һ������
  reg resetSignal_tb;//��������
  reg passwordInputFinishSignal_tb;//������������ź�
  `INPUT_TYPE inputNumber_tb;//����8λ����������

  /* verilator lint_off UNUSEDSIGNAL */
  wire [`PASSWORD_BITS-1:0] display_tb;
  /* verilator lint_off UNUSEDSIGNAL */

  Lock lock (
         .clk(clk_tb),
         .rst_n(rst_n_tb),
         .controlSignal({modeSettingWire_tb, // 3
                         inputNextSignal_tb, // 2 
                         resetSignal_tb, // 1
                         passwordInputFinishSignal_tb}), // 0
         .inputNumber(inputNumber_tb),
         .display(display_tb)
       );//ʵ����Lockģ��

  localparam integer NsPerClk = 1000000;//1ms
  localparam integer NsPerOp = 1000 * NsPerClk;
  always #(NsPerClk / 2) clk_tb = ~clk_tb;//clk_tbÿ1msȡ��


  // ��λ�����������
// `define RANDOM_2_8 ($urandom_range(0, 9)[7:0]*10+$urandom_range(0, 9)[7:0])

  `PASSWORD_TYPE randomPassword;
  `INDEX_TYPE i;


  initial
  begin
    $dumpfile("Lock.vcd");
    $dumpvars(0, tb_Lock);
  end

  initial
  begin
    clk_tb = 0;
    // �����������
    randomPassword = 0;
    // for (i = 0; i < `PASSWORD_LENGTH; i = i + 1)
    fork//fork...join���飬fork...join�����е���䲢��ִ��
      // randomPassword = (randomPassword << 4) + $urandom_range(0, 9)[`PASSWORD_BITS-1:0];
      randomPassword = 24'hCCAA11;
    join

    // ��ʼ��
    fork
      rst_n_tb = 1'b0;
    join
    #NsPerOp;

    // ��ʼִ��
    fork
      rst_n_tb = 1'b1;
    join
    #NsPerOp;

    // ����
    // ��������
    fork
      // inputNumber_tb     = `RANDOM_2_8;
      inputNumber_tb     = 8'hCC;
      inputNextSignal_tb = 1'b1;
    join
    #NsPerOp;

    fork
      // inputNumber_tb     = `RANDOM_2_8;
      inputNumber_tb     = 8'hAA;
      inputNextSignal_tb = 1'b0;
    join
    #NsPerOp;

    fork
      // inputNumber_tb     = `RANDOM_2_8;
      inputNumber_tb     = 8'h11;
      inputNextSignal_tb = 1'b1;
    join
    #NsPerOp;

    fork
      // inputNumber_tb     = `RANDOM_2_8;
      inputNumber_tb     = 8'h11;
      inputNextSignal_tb = 1'b0;
    join
    #NsPerOp;

    // ��������
    fork
      resetSignal_tb = 1'b1;
    join
    #NsPerOp;

    // ��������
    fork
      resetSignal_tb     = 1'b0;
      inputNumber_tb     = randomPassword[23:16];
      inputNextSignal_tb = 1'b1;
    join
    #NsPerOp;

    fork
      inputNumber_tb     = randomPassword[15:8];
      inputNextSignal_tb = 1'b0;
    join
    #NsPerOp;

    fork
      inputNumber_tb     = randomPassword[7:0];
      inputNextSignal_tb = 1'b1;
    join
    #NsPerOp;

    // ����
    fork
      modeSettingWire_tb = 1'b1;
    join
    #NsPerOp;

    // ��������
    fork
      // inputNumber_tb     = `RANDOM_2_8;
      inputNumber_tb     = 8'hCC;
      inputNextSignal_tb = 1'b0;
    join
    #NsPerOp;

    fork
      // inputNumber_tb     = `RANDOM_2_8;
      inputNumber_tb     = 8'hAA;
      inputNextSignal_tb = 1'b1;
    join
    #NsPerOp;

    fork
      // inputNumber_tb     = `RANDOM_2_8;
      inputNumber_tb     = 8'h11;
      inputNextSignal_tb = 1'b0;
    join
    #NsPerOp;

    #NsPerOp;

    // ����������
    fork
      passwordInputFinishSignal_tb = 1'b1;
    join
    #(3.5 * NsPerClk * `CLOCKS_PER_SEC);
    #NsPerOp

     // ��������
     fork
       passwordInputFinishSignal_tb = 1'b0;
       inputNextSignal_tb           = 1'b1;
       inputNumber_tb               = randomPassword[23:16];
     join
     #NsPerOp;

    fork
      inputNextSignal_tb = 1'b0;
      inputNumber_tb     = randomPassword[15:8];
    join
    #NsPerOp;

    fork
      inputNextSignal_tb = 1'b1;
      inputNumber_tb     = randomPassword[7:0];
    join
    #NsPerOp;

    #NsPerOp;

    // �����ȷ����
    fork
      passwordInputFinishSignal_tb = 1'b1;
    join
    #(1.5 * NsPerClk * `CLOCKS_PER_SEC);
    #NsPerOp

     // ���
     fork
       resetSignal_tb = 1'b1;
     join
     #NsPerOp;

    // �ص�����ģʽ
    fork
      modeSettingWire_tb = 1'b0;
    join
    #NsPerOp;

    $finish;
  end

endmodule

/* verilator lint_on BLKSEQ */

`default_nettype wire
